//this is a mux.v file
/* multi
line
comment
*/
module
endmodule
integer 
real

154
5'b10111;
parameter SIZE=32;
session 
book
laptop
verilog
sv
uvm
