module wand_nature(a,b,y);
input a,b;
output y;

assign y=a;
assign y=b;

//assign y=a & b;
//assign y=a | b;
endmodule
