module wor_nature(a,b,y);
input a,b;
output wor y;

//assign y=a;
//assign y=b;

assign y=a & b;
assign y=a | b;

endmodule
