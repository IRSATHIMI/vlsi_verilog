`include "fifo_synch.v"
`include "tb_debug.v"
