`include "mux_4x1.v"
`include "mux_8x1.v"
module tb;



endmodule
