module alu (a,b...., d,e);
  full_adder fa1();
  full_adder fa2();
  multiuplier ma();
endmodule
