`include "sipo_design.v"
module tb;

parameter S_NO_DATA = 3'b001;
parameter S_FETCHING_DATA = 3'b010;
parameter S_WRITE_FIFO = 3'b100;
parameter DEPTH_FIFO = 16;
parameter PCLK_TP = 8;
parameter SCLKTP = 1;

reg sclk_i, pclk_i, rst_i;
reg data_i, valid_i;
wire ready_o;
wire [7:0] data_o;
wire valid_o;
reg ready_i;
integer i ,n;


sipo_design #(.DEPTH_FIFO(DEPTH_FIFO)) dut(sclk_i, pclk_i, rst_i,
data_i, valid_i, ready_o,
data_o, valid_o, ready_i,);

// sclock gen
initial begin
sclk_i =0;
forever #SCLKTP sclk_i = ~sclk_i;
end

// pclock gen
initial begin
pclk_i =0;
forever #PCLK_TP pclk_i = ~pclk_i;
end

initial begin
	// applying reset
	rst_i=1;
	rst_ip();
	repeat (2) @(posedge pclk_i);
	rst_i=0;
	// stimulus;

	for (i=0 ; i<10 ; i=i+1) begin
		@(posedge sclk_i)
		valid_i = 1;
		for(n=0 ; n<=7 ; n=n+1) begin
			@(posedge sclk_i);
			data_i = $random;
			wait (ready_o);
		end
	end
	@(posedge pclk_i);
	valid_i = 0;
	data_i = 0;
		
	#500;
	$finish;
end

task rst_ip();
begin
	data_i = 0;
	valid_i = 0;
	ready_i = 0;
	n=0;
	i=0;
end
endtask

always @(posedge pclk_i) begin
	if(valid_o) ready_i = 1;
	else ready_i = 0;
end
endmodule
